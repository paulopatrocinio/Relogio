--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY display_7segmentos IS
    PORT (
        entrada_display_7segmentos : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		  saida_display_7segmentos : OUT STD_LOGIC_VECTOR (6 DOWNTO 0)
    );
END display_7segmentos;

ARCHITECTURE Behavioral OF display_7segmentos IS
BEGIN
    WITH entrada_display_7segmentos SELECT
        saida_display_7segmentos <= "0000001" WHEN "0000", -- '0'
        "1001111" WHEN "0001", -- '1'
        "0010010" WHEN "0010", -- '2'
        "0000110" WHEN "0011", -- '3'
        "1001100" WHEN "0100", -- '4'
        "0100100" WHEN "0101", -- '5'
        "0100000" WHEN "0110", -- '6'
        "0001111" WHEN "0111", -- '7'
        "0000000" WHEN "1000", -- '8'
        "0000100" WHEN "1001", -- '9'
        "1111111" WHEN OTHERS;
END Behavioral;